module lazy(
    input a,
    input b
);
    
endmodule