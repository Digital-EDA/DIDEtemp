
architecture and_arch of my_entity is
begin
    -- y <= a and b;
end architecture and_arch;

configuration cfg_and_arch of my_entity is
    for and_arch
    end for;
end cfg_and_arch;